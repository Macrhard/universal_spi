module (
    input [79:0]    i_data,
    input []    
);

endmodule // 